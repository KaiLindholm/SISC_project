// ECE:3350 SISC computer project
// finite state machine

`timescale 1ns/100ps



module ctrl (clk, rst_f, opcode, mm, stat, rf_we, alu_op, wb_sel, 
             rb_sel, br_sel, pc_rst, pc_write, pc_sel, ir_load);
  
  input clk, rst_f;
  input [3:0] opcode, mm, stat;
  output reg rf_we, wb_sel, rb_sel, br_sel, pc_rst, pc_write, pc_sel, ir_load;
  output reg [1:0] alu_op;

  // state parameter declarations
  parameter start0 = 0, start1 = 1, fetch = 2, decode = 3, execute = 4, mem = 5, writeback = 6;
   
  // opcode paramenter declarations
  parameter NOOP = 0, LOD = 1, STR = 2, SWP = 3, BRA = 4, BRR = 5, BNE = 6, BNR = 7, ALU_OP = 8, HLT=15;

  // addressing modes
  parameter AM_IMM = 8;

  // state register and next state value
  reg [2:0]  present_state, next_state;

  // Initialize present state to 'start0'.
  initial
    present_state = start0;

  /* Clock procedure that progresses the fsm to the next state on the positive 
     edge of the clock, OR resets the state to 'start1' on the negative edge
     of rst_f. Notice that the computer is reset when rst_f is low, not high. */

  always @(posedge clk, negedge rst_f) begin
    if (rst_f == 1'b0)
      present_state <= start1;
    else
      present_state <= next_state;
  end
  
  /* Combinational procedure that determines the next state of the fsm. */

  always @(present_state, rst_f) begin
    case(present_state)
      start0:
        next_state = start1;
      start1:
	if (rst_f == 1'b0) 
      next_state = start1;
	else
          next_state = fetch;
      fetch:
        next_state = decode;
      decode:
        next_state = execute;
      execute:
        next_state = mem;
      mem:
        next_state = writeback;
      writeback:
        next_state = fetch;
      default:
        next_state = start1;
    endcase
  end
  
  always @(present_state, opcode, mm) begin
    rf_we  = 1'b0;
    wb_sel = 1'b0;
    alu_op = 2'b10;
    rb_sel = 1'b0;
    br_sel = 1'b0; 
    pc_rst = 1'b0; 
    pc_write = 1'b0; 
    pc_sel = 1'b0;
    ir_load = 1'b0;

    case(present_state)
      start1: begin
        pc_rst = 1'b1; 
      end
      fetch: begin
        ir_load = 1'b1; // load the ir with the next instruction 
        pc_sel = 1'b0;  // load PC + 1 
      end

      decode: begin
        if(opcode == BRA) begin 
         if((mm & stat) != 0) begin   // branch taken
              br_sel = 1'b1;    // take branch imm + 0. 
              pc_sel = 1'b1;    // store branch address to pc. 
              pc_write = 1'b1;  // write new value to the pc. 
            end else begin      // the branch is not taken 
              br_sel = 1'b1;    // branch not taken. we want to move ahead in the intrusctions
              //pc_sel = 1'b0;    // PC + 1 
              pc_write = 1'b1;  // write the new value to PC 
            end 
        end else if(opcode == BRR) begin 
          if((mm & stat) != 0) begin    // branch taken 
                  pc_sel = 1'b1; // save the branch address to pc 
                  br_sel = 1'b1; // branch address is imm + PC + 1
                  pc_write = 1'b1; // write new value to the pc. 
          end else begin  // the branch is not taken 
                  //pc_sel = 1'b0; // write PC + 1 to the pc 
                  br_sel = 1'b1; // branch not taken. we want to move ahead in the intrusctions 
                  pc_write = 1'b1;  // write the new value to PC 
          end
        end else if(opcode == BNE) begin 
          if((mm & stat) == 0) begin    //  branch is not taken 
                pc_sel = 1'b0; // write PC + 1 to the pc 
                br_sel = 1'b1; // branch not taken. we want to move ahead in the intrusctions 
                pc_write = 1'b1;  // write the new value to PC 
              end else begin  // the branch is taken 
                pc_sel = 1'b1; // save the branch address to pc 
                br_sel = 1'b1; // absolute branching. 
                pc_write = 1'b1; // write new value to the pc. 
              end
        end else if(opcode == BNR) begin 
          if((4'b0010 & stat) == 0) begin    //  branch is not taken 
                pc_sel = 1'b0; // next instruciton 
                br_sel = 1'b1; // add pc + 1 to 0. 
                pc_write = 1'b1;  // write the new value to PC 
              end else begin  // the branch is taken 
                pc_sel = 1'b1; // save the branch address to pc 
                br_sel = 1'b0; // relative branching. 
                pc_write = 1'b1; // write new value to the pc. 
              end
        end else begin 
          pc_sel = 1'b0; // next instruction is taken 
              br_sel = 1'b1; 
              pc_write = 1'b1; 
        end 
      end

      execute: begin
        if ((opcode == ALU_OP) && (mm == AM_IMM))
          alu_op = 2'b01;
        else
          alu_op = 2'b00;
      end

      mem: begin
        if ((opcode == ALU_OP) && (mm == AM_IMM))
          alu_op = 2'b11;
        else
          alu_op = 2'b10;
      end

      writeback: begin
        if (opcode == ALU_OP)
          rf_we = 1'b1;  
      end

      default: begin
        rf_we  = 1'b0;
        wb_sel = 1'b0;
        alu_op = 2'b10;
        rb_sel = 1'b0;
        br_sel = 1'b0; 
        pc_rst = 1'b0; 
        pc_write = 1'b0; 
        pc_sel = 1'b0;
        ir_load = 1'b0;
      end
    endcase
  end

// Halt on HLT instruction  
  always @(opcode)
  begin
    if (opcode == HLT)
    begin 
      #5 $display ("Halt."); //Delay 5 ns so $monitor will print the halt instruction
      $stop;
    end
  end
    
  
endmodule
